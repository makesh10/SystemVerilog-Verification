interface inter();
  logic clk;
  logic rst;
  logic counter;
  logic [6:0]count;
endinterface
